module controlunit (
    input logic [31:0] instruction,
    input logic eq,
    output logic regwrite, alusrc, pcsrc, memwrite, resultsrc,
    output logic [2:0] aluctrl, immsrc, addrmode
);

  
endmodule
