module name #(
    parameters D_WIDTH
) (
    input 
);
    
endmodule