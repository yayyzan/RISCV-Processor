module controlunit (
    input logic [31:0] instruction,
    input logic eq,
    output logic regwrite,
    output logic [2:0] aluctrl,
    output logic alusrc,
    output logic pcsrc,
    output logic [2:0] immsrc,
    output logic memwrite,
    output logic [2:0] addrmode,
    output logic resultsrc
);


endmodule
